module Program_Counter_tb;

