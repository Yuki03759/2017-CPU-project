module barrel_tb;

