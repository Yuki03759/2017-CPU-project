module example1