module example_fulladder();


