module XOR_Tree